

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO system_top_dft 
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.383 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.84223 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.23232 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 23.756 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 114.459 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 581.907 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2816.37 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 2.383 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4622 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.26022 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.584 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.4314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 14.736 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 71.0726 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 8.996 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 43.4632 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 443.539 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 2150.82 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA67 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 2.005 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.64405 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.042 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.20442 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.192 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7859 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 152.038 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 741.483 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[0]
  PIN SO[2] 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 1.424 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.84944 LAYER METAL3 ;
  END SO[2]
  PIN SO[0] 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 0.194 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL3 ;
  END SO[0]
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.455 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.18855 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.534 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.57094 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.635889 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 3.14155 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.141 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.67821 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.561 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.70081 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.644704 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 3.18396 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END UART_CLK
  PIN RST 
    ANTENNAPARTIALMETALAREA 3.452 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6041 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.367 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.15007 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 24.8405 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 126.846 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END RST
  PIN RX_IN 
    ANTENNAPARTIALMETALAREA 1.352 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 6.50312 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.88 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.43 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7761 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 13.5548 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 65.7653 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA34 ;
  END RX_IN
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.237 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.13997 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.02116 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 11.957 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 57.7056 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.247 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 112.874 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 545.181 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.78775 LAYER VIA56 ;
  END SE
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.419 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.01539 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.41558 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.421706 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2.11133 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 0.223 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.07263 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 12.768 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.6065 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 232.076 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1122.45 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.48343 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 3.649 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5517 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 24.7675 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 117.37 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.205698 LAYER VIA23 ;
  END test_mode
  PIN TX_OUT 
    ANTENNAPARTIALMETALAREA 0.86 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1366 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.26022 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.537 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 7.766 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 37.5469 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 153.878 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 749.512 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END TX_OUT
  PIN PAR_ERR 
    ANTENNAPARTIALMETALAREA 0.86 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.1366 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNADIFFAREA 0.6 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 6.102 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7354 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5239 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 40.3556 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 197.006 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.63368 LAYER VIA45 ;
  END PAR_ERR
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 29.609 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 142.997 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 421.781 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2036.99 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.514245 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 5.962 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8696 LAYER METAL4 ;
    ANTENNAGATEAREA 0.1404 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 464.245 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 2242.61 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.54274 LAYER VIA45 ;
  END SO[1]
  PIN STP_ERR 
    ANTENNAPARTIALMETALAREA 2.089 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4329 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 31.9188 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 156.706 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 1.54274 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 29.629 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 143.093 LAYER METAL3 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 453.984 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2195.06 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.05698 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 5.962 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 28.8696 LAYER METAL4 ;
    ANTENNAGATEAREA 0.1404 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 496.449 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 2400.69 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.05698 LAYER VIA45 ;
  END STP_ERR
END system_top_dft

END LIBRARY
