module UART_RX #(parameter width=8)(
input wire CLK,RST,  
input wire RX_IN,
input wire [5:0] PRESCALE,
input wire PAR_TYP,
input wire PAR_EN,
output wire DATA_VALID,
output wire [width-1:0] P_DATA,  
output wire PAR_ERR,
output wire STP_ERR
);

wire ENABLE,DATA_SAMP_EN,SAMPLED_BIT,PAR_CHK_EN,STRT_CHK_EN,STRT_GLITCH;
wire STP_CHK_EN,DESER_EN;
wire [3:0] BIT_CNT;
wire [4:0] EDGE_CNT;

FSM F (
.RX_IN(RX_IN),
.CLK(CLK),
.RST(RST),
.PAR_EN(PAR_EN),
.BIT_CNT(BIT_CNT),
.PAR_ERR(PAR_ERR),
.STRT_GLITCH(STRT_GLITCH),
.STP_ERR(STP_ERR),
.ENABLE(ENABLE),
.DATA_SAMP_EN(DATA_SAMP_EN),
.DESER_EN(DESER_EN),
.DATA_VALID(DATA_VALID),
.PAR_CHK_EN(PAR_CHK_EN),
.STRT_CHK_EN(STRT_CHK_EN),
.STP_CHK_EN(STP_CHK_EN),
.PRESCALE(PRESCALE),
.EDGE_CNT(EDGE_CNT)
);

data_sampling D0 (
.RX_IN(RX_IN),
.CLK(CLK),
.RST(RST),
.PRESCALE(PRESCALE),
.DATA_SAMP_EN(DATA_SAMP_EN),
.EDGE_CNT(EDGE_CNT),
.SAMPLED_BIT(SAMPLED_BIT)
);

deserializer D1 (
.CLK(CLK),
.RST(RST),
.SAMPLED_BIT(SAMPLED_BIT),
.DESER_EN(DESER_EN),
.P_DATA(P_DATA)
);

edge_bit_counter E(
.CLK(CLK),
.RST(RST),
.PAR_EN(PAR_EN),
.ENABLE(ENABLE),
.PRESCALE(PRESCALE),
.EDGE_CNT(EDGE_CNT),
.BIT_CNT(BIT_CNT)
);

PARITY_CHECK P(
.CLK(CLK),
.RST(RST),
.SAMPLED_BIT(SAMPLED_BIT),
.P_DATA(P_DATA),
.PAR_CHK_EN(PAR_CHK_EN),
.PAR_TYP(PAR_TYP),
.PAR_ERR(PAR_ERR)
);

STRT_CHECK S0(
.CLK(CLK),
.RST(RST),
.SAMPLED_BIT(SAMPLED_BIT),
.STRT_CHK_EN(STRT_CHK_EN),
.STRT_GLITCH(STRT_GLITCH)
);

STOP_CHECK S1 (
.CLK(CLK),
.RST(RST),
.SAMPLED_BIT(SAMPLED_BIT),
.STP_CHK_EN(STP_CHK_EN),
.STP_ERR(STP_ERR)
);

endmodule